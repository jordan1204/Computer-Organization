
module INSTRUCTION_FETCH(
	clk,
	rst,
	jump,
	branch,
	jump_addr,
	branch_addr,

	PC,
	IR
);

input clk, rst, jump, branch;
input [31:0] jump_addr, branch_addr;

output reg 	[31:0] PC;
output reg 	[31:0] IR;

reg [31:0] instruction [127:0];
//output instruction
always @(posedge clk or posedge rst)
begin
	if(rst) begin
		IR <= 32'd0;
	    instruction[0 ] <= 32'b100011_00000_00011_00000_00000_000000;  //Lw mem0 to r3
        instruction[1 ] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[2 ] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[3 ] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[4 ] <= 32'b000000_00011_00000_01001_00000_100000;    //copy r3 to t1 (add)
        instruction[5 ] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[6 ] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[7 ] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)        
        instruction[8 ] <= 32'b000000_00011_00000_01111_00000_100000;    //copy r3 to t7 (add)
        instruction[9 ] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[10] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[11] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)    
        instruction[12] <= 32'b000000_01001_00001_01001_00000_100010;    //sub t1 1       //next1
        instruction[13] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[14] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[15] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)        
        instruction[16] <= 32'b000100_01001_00010_0000000000110011;    //beq t1, $2, 40 
        instruction[17] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[18] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[19] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[20] <= 32'b000000_00000_00010_01011_00000_100000;    //addi t3 2      
        instruction[21] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[22] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[23] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)    
        instruction[24] <= 32'b000000_00000_01001_01110_00000_100000;    //add t6 t1 0    //sub 1
        instruction[25] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[26] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[27] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)    
        instruction[28] <= 32'b000000_01110_01011_01110_00000_100010;    //sub t6 t6 t3    //div 1
        instruction[29] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[30] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[31] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[32] <= 32'b000100_01110_00000_1111111111101010;    //beq t6, 0, -22
        instruction[33] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[34] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[35] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[36] <= 32'b000000_01110_01011_10000_00000_101010;    //slt t8, t6, t3              t8 = 1
        instruction[37] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[38] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[39] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[40] <= 32'b000100_10000_00000_11111_11111_110010;    //beq t8, 0, -14
        instruction[41] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[42] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[43] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[44] <= 32'b000000_01011_00001_01011_00000_100000;    //add t3 t3 1 (add)
        instruction[45] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[46] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[47] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[48] <= 32'b000000_01011_01011_01100_00000_100000;    //add t4 t3 t3 (add)
        instruction[49] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[50] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[51] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[52] <= 32'b000100_01001_01100_11111_11111_010111;    //beq t4, t1, -40
        instruction[53] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[54] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[55] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[56] <= 32'b000000_01100_01001_01101_00000_101010;    //slt t4, t1, t5              t5 = 1
        instruction[57] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[58] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[59] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[60] <= 32'b000100_01101_00000_00000_00000_000111;    //beq t5, 0, next 2 
        instruction[61] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[62] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[63] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[64] <= 32'b000010_00000_00000_00000_00000_010111;    //j 23                // j sub
        instruction[65] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[66] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[67] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[68] <= 32'b000000_01111_00001_01111_00000_100000;    //add t7 1           //next2
        instruction[69] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[70] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[71] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)        
        instruction[72] <= 32'b000000_00000_00010_01011_00000_100000;    //add t3 0  2      
        instruction[73] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[74] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[75] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)    
        instruction[76] <= 32'b000000_00000_01111_01110_00000_100000;    //add t6 t7 0    //add 1
        instruction[77] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[78] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[79] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)    
        instruction[80] <= 32'b000000_01110_01011_01110_00000_100010;    //sub t6 t6 t3    //div 2
        instruction[81] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[82] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[83] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[84] <= 32'b000100_01110_00000_1111111111101111;    //beq t6, 0, next2 
        instruction[85] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[86] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[87] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[88] <= 32'b000000_01110_01011_10000_00000_101010;    //slt t8, t6, t3              t8 = 1
        instruction[89] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[90] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[91] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[92] <= 32'b000100_10000_00000_1111111111110011;    //beq t8, 0, div2
        instruction[93] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[94] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[95] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[96] <= 32'b000000_01011_00001_01011_00000_100000;    //add t3 t3 1 (add)
        instruction[97] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[98] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[99] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[100] <= 32'b000000_01011_01011_01100_00000_100000;    //add t4 t3 t3 (add)
        instruction[101] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[102] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[103] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[104] <= 32'b000100_01100_01111_1111111111101100;    //beq $t4,$t7,next2
        instruction[105] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[106] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[107] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[108] <= 32'b000000_01100_01111_01101_00000_101010;    //slt $t5,$t4,$t7
        instruction[109] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[110] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[111] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[112] <= 32'b000100_01101_00000_00000_00000_000111;    //beq t5, 0, 7
        instruction[113] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[114] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[115] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[116] <= 32'b000010_00000_00000_00000_00001_001011;    //j add1
        instruction[117] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[118] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[119] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[120] <= 32'b101011_00000_01001_0000000000000010;    //SW $1, 3                
        instruction[121] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[122] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[123] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[124] <= 32'b101011_00000_01111_0000000000000011;    //SW $7, 4               
        instruction[125] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[126] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[127] <= 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
	end
	else begin
		if(PC[10:2]<=8'd127) 
		  IR <= instruction[PC[10:2]]; //(0, 4, 8, ...) => (0, 1, 2, ...)
		//else
		  //IR <= IR;
	end
end

// output program counter
always @(posedge clk or posedge rst)
begin
	if(rst)
		PC <= 32'd0;
	else begin
	   if(PC[10:2]<8'd127) 
	       PC <= (branch) ? branch_addr : ( (jump) ? jump_addr : (PC+4)) ;
	   //else
	       //PC <= PC;
	end
end

endmodule